module PaletasLimites(input [11:0] contador,output reg[10:0] saidaYMax,saidaYm);
always @ (contador)
begin
case(contador)
0:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
1:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
2:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
3:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
4:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
5:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
6:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
7:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
8:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
9:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
10:
    begin
        saidaYMax<=95;
        saidaYm<=5;
    end
11:
    begin
        saidaYMax<=96;
        saidaYm<=6;
    end
12:
    begin
        saidaYMax<=96;
        saidaYm<=6;
    end
13:
    begin
        saidaYMax<=96;
        saidaYm<=6;
    end
14:
    begin
        saidaYMax<=96;
        saidaYm<=6;
    end
15:
    begin
        saidaYMax<=96;
        saidaYm<=6;
    end
16:
    begin
        saidaYMax<=96;
        saidaYm<=6;
    end
17:
    begin
        saidaYMax<=96;
        saidaYm<=6;
    end
18:
    begin
        saidaYMax<=96;
        saidaYm<=6;
    end
19:
    begin
        saidaYMax<=96;
        saidaYm<=6;
    end
20:
    begin
        saidaYMax<=96;
        saidaYm<=6;
    end
21:
    begin
        saidaYMax<=97;
        saidaYm<=7;
    end
22:
    begin
        saidaYMax<=97;
        saidaYm<=7;
    end
23:
    begin
        saidaYMax<=97;
        saidaYm<=7;
    end
24:
    begin
        saidaYMax<=97;
        saidaYm<=7;
    end
25:
    begin
        saidaYMax<=97;
        saidaYm<=7;
    end
26:
    begin
        saidaYMax<=97;
        saidaYm<=7;
    end
27:
    begin
        saidaYMax<=97;
        saidaYm<=7;
    end
28:
    begin
        saidaYMax<=97;
        saidaYm<=7;
    end
29:
    begin
        saidaYMax<=97;
        saidaYm<=7;
    end
30:
    begin
        saidaYMax<=97;
        saidaYm<=7;
    end
31:
    begin
        saidaYMax<=98;
        saidaYm<=8;
    end
32:
    begin
        saidaYMax<=98;
        saidaYm<=8;
    end
33:
    begin
        saidaYMax<=98;
        saidaYm<=8;
    end
34:
    begin
        saidaYMax<=98;
        saidaYm<=8;
    end
35:
    begin
        saidaYMax<=98;
        saidaYm<=8;
    end
36:
    begin
        saidaYMax<=98;
        saidaYm<=8;
    end
37:
    begin
        saidaYMax<=98;
        saidaYm<=8;
    end
38:
    begin
        saidaYMax<=98;
        saidaYm<=8;
    end
39:
    begin
        saidaYMax<=98;
        saidaYm<=8;
    end
40:
    begin
        saidaYMax<=98;
        saidaYm<=8;
    end
41:
    begin
        saidaYMax<=99;
        saidaYm<=9;
    end
42:
    begin
        saidaYMax<=99;
        saidaYm<=9;
    end
43:
    begin
        saidaYMax<=99;
        saidaYm<=9;
    end
44:
    begin
        saidaYMax<=99;
        saidaYm<=9;
    end
45:
    begin
        saidaYMax<=99;
        saidaYm<=9;
    end
46:
    begin
        saidaYMax<=99;
        saidaYm<=9;
    end
47:
    begin
        saidaYMax<=99;
        saidaYm<=9;
    end
48:
    begin
        saidaYMax<=99;
        saidaYm<=9;
    end
49:
    begin
        saidaYMax<=99;
        saidaYm<=9;
    end
50:
    begin
        saidaYMax<=99;
        saidaYm<=9;
    end
51:
    begin
        saidaYMax<=100;
        saidaYm<=10;
    end
52:
    begin
        saidaYMax<=100;
        saidaYm<=10;
    end
53:
    begin
        saidaYMax<=100;
        saidaYm<=10;
    end
54:
    begin
        saidaYMax<=100;
        saidaYm<=10;
    end
55:
    begin
        saidaYMax<=100;
        saidaYm<=10;
    end
56:
    begin
        saidaYMax<=100;
        saidaYm<=10;
    end
57:
    begin
        saidaYMax<=100;
        saidaYm<=10;
    end
58:
    begin
        saidaYMax<=100;
        saidaYm<=10;
    end
59:
    begin
        saidaYMax<=100;
        saidaYm<=10;
    end
60:
    begin
        saidaYMax<=100;
        saidaYm<=10;
    end
61:
    begin
        saidaYMax<=101;
        saidaYm<=11;
    end
62:
    begin
        saidaYMax<=101;
        saidaYm<=11;
    end
63:
    begin
        saidaYMax<=101;
        saidaYm<=11;
    end
64:
    begin
        saidaYMax<=101;
        saidaYm<=11;
    end
65:
    begin
        saidaYMax<=101;
        saidaYm<=11;
    end
66:
    begin
        saidaYMax<=101;
        saidaYm<=11;
    end
67:
    begin
        saidaYMax<=101;
        saidaYm<=11;
    end
68:
    begin
        saidaYMax<=101;
        saidaYm<=11;
    end
69:
    begin
        saidaYMax<=101;
        saidaYm<=11;
    end
70:
    begin
        saidaYMax<=101;
        saidaYm<=11;
    end
71:
    begin
        saidaYMax<=102;
        saidaYm<=12;
    end
72:
    begin
        saidaYMax<=102;
        saidaYm<=12;
    end
73:
    begin
        saidaYMax<=102;
        saidaYm<=12;
    end
74:
    begin
        saidaYMax<=102;
        saidaYm<=12;
    end
75:
    begin
        saidaYMax<=102;
        saidaYm<=12;
    end
76:
    begin
        saidaYMax<=102;
        saidaYm<=12;
    end
77:
    begin
        saidaYMax<=102;
        saidaYm<=12;
    end
78:
    begin
        saidaYMax<=102;
        saidaYm<=12;
    end
79:
    begin
        saidaYMax<=102;
        saidaYm<=12;
    end
80:
    begin
        saidaYMax<=102;
        saidaYm<=12;
    end
81:
    begin
        saidaYMax<=103;
        saidaYm<=13;
    end
82:
    begin
        saidaYMax<=103;
        saidaYm<=13;
    end
83:
    begin
        saidaYMax<=103;
        saidaYm<=13;
    end
84:
    begin
        saidaYMax<=103;
        saidaYm<=13;
    end
85:
    begin
        saidaYMax<=103;
        saidaYm<=13;
    end
86:
    begin
        saidaYMax<=103;
        saidaYm<=13;
    end
87:
    begin
        saidaYMax<=103;
        saidaYm<=13;
    end
88:
    begin
        saidaYMax<=103;
        saidaYm<=13;
    end
89:
    begin
        saidaYMax<=103;
        saidaYm<=13;
    end
90:
    begin
        saidaYMax<=103;
        saidaYm<=13;
    end
91:
    begin
        saidaYMax<=104;
        saidaYm<=14;
    end
92:
    begin
        saidaYMax<=104;
        saidaYm<=14;
    end
93:
    begin
        saidaYMax<=104;
        saidaYm<=14;
    end
94:
    begin
        saidaYMax<=104;
        saidaYm<=14;
    end
95:
    begin
        saidaYMax<=104;
        saidaYm<=14;
    end
96:
    begin
        saidaYMax<=104;
        saidaYm<=14;
    end
97:
    begin
        saidaYMax<=104;
        saidaYm<=14;
    end
98:
    begin
        saidaYMax<=104;
        saidaYm<=14;
    end
99:
    begin
        saidaYMax<=104;
        saidaYm<=14;
    end
100:
    begin
        saidaYMax<=104;
        saidaYm<=14;
    end
101:
    begin
        saidaYMax<=105;
        saidaYm<=15;
    end
102:
    begin
        saidaYMax<=105;
        saidaYm<=15;
    end
103:
    begin
        saidaYMax<=105;
        saidaYm<=15;
    end
104:
    begin
        saidaYMax<=105;
        saidaYm<=15;
    end
105:
    begin
        saidaYMax<=105;
        saidaYm<=15;
    end
106:
    begin
        saidaYMax<=105;
        saidaYm<=15;
    end
107:
    begin
        saidaYMax<=105;
        saidaYm<=15;
    end
108:
    begin
        saidaYMax<=105;
        saidaYm<=15;
    end
109:
    begin
        saidaYMax<=105;
        saidaYm<=15;
    end
110:
    begin
        saidaYMax<=105;
        saidaYm<=15;
    end
111:
    begin
        saidaYMax<=106;
        saidaYm<=16;
    end
112:
    begin
        saidaYMax<=106;
        saidaYm<=16;
    end
113:
    begin
        saidaYMax<=106;
        saidaYm<=16;
    end
114:
    begin
        saidaYMax<=106;
        saidaYm<=16;
    end
115:
    begin
        saidaYMax<=106;
        saidaYm<=16;
    end
116:
    begin
        saidaYMax<=106;
        saidaYm<=16;
    end
117:
    begin
        saidaYMax<=106;
        saidaYm<=16;
    end
118:
    begin
        saidaYMax<=106;
        saidaYm<=16;
    end
119:
    begin
        saidaYMax<=106;
        saidaYm<=16;
    end
120:
    begin
        saidaYMax<=106;
        saidaYm<=16;
    end
121:
    begin
        saidaYMax<=107;
        saidaYm<=17;
    end
122:
    begin
        saidaYMax<=107;
        saidaYm<=17;
    end
123:
    begin
        saidaYMax<=107;
        saidaYm<=17;
    end
124:
    begin
        saidaYMax<=107;
        saidaYm<=17;
    end
125:
    begin
        saidaYMax<=107;
        saidaYm<=17;
    end
126:
    begin
        saidaYMax<=107;
        saidaYm<=17;
    end
127:
    begin
        saidaYMax<=107;
        saidaYm<=17;
    end
128:
    begin
        saidaYMax<=107;
        saidaYm<=17;
    end
129:
    begin
        saidaYMax<=107;
        saidaYm<=17;
    end
130:
    begin
        saidaYMax<=107;
        saidaYm<=17;
    end
131:
    begin
        saidaYMax<=108;
        saidaYm<=18;
    end
132:
    begin
        saidaYMax<=108;
        saidaYm<=18;
    end
133:
    begin
        saidaYMax<=108;
        saidaYm<=18;
    end
134:
    begin
        saidaYMax<=108;
        saidaYm<=18;
    end
135:
    begin
        saidaYMax<=108;
        saidaYm<=18;
    end
136:
    begin
        saidaYMax<=108;
        saidaYm<=18;
    end
137:
    begin
        saidaYMax<=108;
        saidaYm<=18;
    end
138:
    begin
        saidaYMax<=108;
        saidaYm<=18;
    end
139:
    begin
        saidaYMax<=108;
        saidaYm<=18;
    end
140:
    begin
        saidaYMax<=108;
        saidaYm<=18;
    end
141:
    begin
        saidaYMax<=109;
        saidaYm<=19;
    end
142:
    begin
        saidaYMax<=109;
        saidaYm<=19;
    end
143:
    begin
        saidaYMax<=109;
        saidaYm<=19;
    end
144:
    begin
        saidaYMax<=109;
        saidaYm<=19;
    end
145:
    begin
        saidaYMax<=109;
        saidaYm<=19;
    end
146:
    begin
        saidaYMax<=109;
        saidaYm<=19;
    end
147:
    begin
        saidaYMax<=109;
        saidaYm<=19;
    end
148:
    begin
        saidaYMax<=109;
        saidaYm<=19;
    end
149:
    begin
        saidaYMax<=109;
        saidaYm<=19;
    end
150:
    begin
        saidaYMax<=109;
        saidaYm<=19;
    end
151:
    begin
        saidaYMax<=110;
        saidaYm<=20;
    end
152:
    begin
        saidaYMax<=110;
        saidaYm<=20;
    end
153:
    begin
        saidaYMax<=110;
        saidaYm<=20;
    end
154:
    begin
        saidaYMax<=110;
        saidaYm<=20;
    end
155:
    begin
        saidaYMax<=110;
        saidaYm<=20;
    end
156:
    begin
        saidaYMax<=110;
        saidaYm<=20;
    end
157:
    begin
        saidaYMax<=110;
        saidaYm<=20;
    end
158:
    begin
        saidaYMax<=110;
        saidaYm<=20;
    end
159:
    begin
        saidaYMax<=110;
        saidaYm<=20;
    end
160:
    begin
        saidaYMax<=110;
        saidaYm<=20;
    end
161:
    begin
        saidaYMax<=111;
        saidaYm<=21;
    end
162:
    begin
        saidaYMax<=111;
        saidaYm<=21;
    end
163:
    begin
        saidaYMax<=111;
        saidaYm<=21;
    end
164:
    begin
        saidaYMax<=111;
        saidaYm<=21;
    end
165:
    begin
        saidaYMax<=111;
        saidaYm<=21;
    end
166:
    begin
        saidaYMax<=111;
        saidaYm<=21;
    end
167:
    begin
        saidaYMax<=111;
        saidaYm<=21;
    end
168:
    begin
        saidaYMax<=111;
        saidaYm<=21;
    end
169:
    begin
        saidaYMax<=111;
        saidaYm<=21;
    end
170:
    begin
        saidaYMax<=111;
        saidaYm<=21;
    end
171:
    begin
        saidaYMax<=112;
        saidaYm<=22;
    end
172:
    begin
        saidaYMax<=112;
        saidaYm<=22;
    end
173:
    begin
        saidaYMax<=112;
        saidaYm<=22;
    end
174:
    begin
        saidaYMax<=112;
        saidaYm<=22;
    end
175:
    begin
        saidaYMax<=112;
        saidaYm<=22;
    end
176:
    begin
        saidaYMax<=112;
        saidaYm<=22;
    end
177:
    begin
        saidaYMax<=112;
        saidaYm<=22;
    end
178:
    begin
        saidaYMax<=112;
        saidaYm<=22;
    end
179:
    begin
        saidaYMax<=112;
        saidaYm<=22;
    end
180:
    begin
        saidaYMax<=112;
        saidaYm<=22;
    end
181:
    begin
        saidaYMax<=113;
        saidaYm<=23;
    end
182:
    begin
        saidaYMax<=113;
        saidaYm<=23;
    end
183:
    begin
        saidaYMax<=113;
        saidaYm<=23;
    end
184:
    begin
        saidaYMax<=113;
        saidaYm<=23;
    end
185:
    begin
        saidaYMax<=113;
        saidaYm<=23;
    end
186:
    begin
        saidaYMax<=113;
        saidaYm<=23;
    end
187:
    begin
        saidaYMax<=113;
        saidaYm<=23;
    end
188:
    begin
        saidaYMax<=113;
        saidaYm<=23;
    end
189:
    begin
        saidaYMax<=113;
        saidaYm<=23;
    end
190:
    begin
        saidaYMax<=113;
        saidaYm<=23;
    end
191:
    begin
        saidaYMax<=114;
        saidaYm<=24;
    end
192:
    begin
        saidaYMax<=114;
        saidaYm<=24;
    end
193:
    begin
        saidaYMax<=114;
        saidaYm<=24;
    end
194:
    begin
        saidaYMax<=114;
        saidaYm<=24;
    end
195:
    begin
        saidaYMax<=114;
        saidaYm<=24;
    end
196:
    begin
        saidaYMax<=114;
        saidaYm<=24;
    end
197:
    begin
        saidaYMax<=114;
        saidaYm<=24;
    end
198:
    begin
        saidaYMax<=114;
        saidaYm<=24;
    end
199:
    begin
        saidaYMax<=114;
        saidaYm<=24;
    end
200:
    begin
        saidaYMax<=114;
        saidaYm<=24;
    end
201:
    begin
        saidaYMax<=115;
        saidaYm<=25;
    end
202:
    begin
        saidaYMax<=115;
        saidaYm<=25;
    end
203:
    begin
        saidaYMax<=115;
        saidaYm<=25;
    end
204:
    begin
        saidaYMax<=115;
        saidaYm<=25;
    end
205:
    begin
        saidaYMax<=115;
        saidaYm<=25;
    end
206:
    begin
        saidaYMax<=115;
        saidaYm<=25;
    end
207:
    begin
        saidaYMax<=115;
        saidaYm<=25;
    end
208:
    begin
        saidaYMax<=115;
        saidaYm<=25;
    end
209:
    begin
        saidaYMax<=115;
        saidaYm<=25;
    end
210:
    begin
        saidaYMax<=115;
        saidaYm<=25;
    end
211:
    begin
        saidaYMax<=116;
        saidaYm<=26;
    end
212:
    begin
        saidaYMax<=116;
        saidaYm<=26;
    end
213:
    begin
        saidaYMax<=116;
        saidaYm<=26;
    end
214:
    begin
        saidaYMax<=116;
        saidaYm<=26;
    end
215:
    begin
        saidaYMax<=116;
        saidaYm<=26;
    end
216:
    begin
        saidaYMax<=116;
        saidaYm<=26;
    end
217:
    begin
        saidaYMax<=116;
        saidaYm<=26;
    end
218:
    begin
        saidaYMax<=116;
        saidaYm<=26;
    end
219:
    begin
        saidaYMax<=116;
        saidaYm<=26;
    end
220:
    begin
        saidaYMax<=116;
        saidaYm<=26;
    end
221:
    begin
        saidaYMax<=117;
        saidaYm<=27;
    end
222:
    begin
        saidaYMax<=117;
        saidaYm<=27;
    end
223:
    begin
        saidaYMax<=117;
        saidaYm<=27;
    end
224:
    begin
        saidaYMax<=117;
        saidaYm<=27;
    end
225:
    begin
        saidaYMax<=117;
        saidaYm<=27;
    end
226:
    begin
        saidaYMax<=117;
        saidaYm<=27;
    end
227:
    begin
        saidaYMax<=117;
        saidaYm<=27;
    end
228:
    begin
        saidaYMax<=117;
        saidaYm<=27;
    end
229:
    begin
        saidaYMax<=117;
        saidaYm<=27;
    end
230:
    begin
        saidaYMax<=117;
        saidaYm<=27;
    end
231:
    begin
        saidaYMax<=118;
        saidaYm<=28;
    end
232:
    begin
        saidaYMax<=118;
        saidaYm<=28;
    end
233:
    begin
        saidaYMax<=118;
        saidaYm<=28;
    end
234:
    begin
        saidaYMax<=118;
        saidaYm<=28;
    end
235:
    begin
        saidaYMax<=118;
        saidaYm<=28;
    end
236:
    begin
        saidaYMax<=118;
        saidaYm<=28;
    end
237:
    begin
        saidaYMax<=118;
        saidaYm<=28;
    end
238:
    begin
        saidaYMax<=118;
        saidaYm<=28;
    end
239:
    begin
        saidaYMax<=118;
        saidaYm<=28;
    end
240:
    begin
        saidaYMax<=118;
        saidaYm<=28;
    end
241:
    begin
        saidaYMax<=119;
        saidaYm<=29;
    end
242:
    begin
        saidaYMax<=119;
        saidaYm<=29;
    end
243:
    begin
        saidaYMax<=119;
        saidaYm<=29;
    end
244:
    begin
        saidaYMax<=119;
        saidaYm<=29;
    end
245:
    begin
        saidaYMax<=119;
        saidaYm<=29;
    end
246:
    begin
        saidaYMax<=119;
        saidaYm<=29;
    end
247:
    begin
        saidaYMax<=119;
        saidaYm<=29;
    end
248:
    begin
        saidaYMax<=119;
        saidaYm<=29;
    end
249:
    begin
        saidaYMax<=119;
        saidaYm<=29;
    end
250:
    begin
        saidaYMax<=119;
        saidaYm<=29;
    end
251:
    begin
        saidaYMax<=120;
        saidaYm<=30;
    end
252:
    begin
        saidaYMax<=120;
        saidaYm<=30;
    end
253:
    begin
        saidaYMax<=120;
        saidaYm<=30;
    end
254:
    begin
        saidaYMax<=120;
        saidaYm<=30;
    end
255:
    begin
        saidaYMax<=120;
        saidaYm<=30;
    end
256:
    begin
        saidaYMax<=120;
        saidaYm<=30;
    end
257:
    begin
        saidaYMax<=120;
        saidaYm<=30;
    end
258:
    begin
        saidaYMax<=120;
        saidaYm<=30;
    end
259:
    begin
        saidaYMax<=120;
        saidaYm<=30;
    end
260:
    begin
        saidaYMax<=120;
        saidaYm<=30;
    end
261:
    begin
        saidaYMax<=121;
        saidaYm<=31;
    end
262:
    begin
        saidaYMax<=121;
        saidaYm<=31;
    end
263:
    begin
        saidaYMax<=121;
        saidaYm<=31;
    end
264:
    begin
        saidaYMax<=121;
        saidaYm<=31;
    end
265:
    begin
        saidaYMax<=121;
        saidaYm<=31;
    end
266:
    begin
        saidaYMax<=121;
        saidaYm<=31;
    end
267:
    begin
        saidaYMax<=121;
        saidaYm<=31;
    end
268:
    begin
        saidaYMax<=121;
        saidaYm<=31;
    end
269:
    begin
        saidaYMax<=121;
        saidaYm<=31;
    end
270:
    begin
        saidaYMax<=121;
        saidaYm<=31;
    end
271:
    begin
        saidaYMax<=122;
        saidaYm<=32;
    end
272:
    begin
        saidaYMax<=122;
        saidaYm<=32;
    end
273:
    begin
        saidaYMax<=122;
        saidaYm<=32;
    end
274:
    begin
        saidaYMax<=122;
        saidaYm<=32;
    end
275:
    begin
        saidaYMax<=122;
        saidaYm<=32;
    end
276:
    begin
        saidaYMax<=122;
        saidaYm<=32;
    end
277:
    begin
        saidaYMax<=122;
        saidaYm<=32;
    end
278:
    begin
        saidaYMax<=122;
        saidaYm<=32;
    end
279:
    begin
        saidaYMax<=122;
        saidaYm<=32;
    end
280:
    begin
        saidaYMax<=122;
        saidaYm<=32;
    end
281:
    begin
        saidaYMax<=123;
        saidaYm<=33;
    end
282:
    begin
        saidaYMax<=123;
        saidaYm<=33;
    end
283:
    begin
        saidaYMax<=123;
        saidaYm<=33;
    end
284:
    begin
        saidaYMax<=123;
        saidaYm<=33;
    end
285:
    begin
        saidaYMax<=123;
        saidaYm<=33;
    end
286:
    begin
        saidaYMax<=123;
        saidaYm<=33;
    end
287:
    begin
        saidaYMax<=123;
        saidaYm<=33;
    end
288:
    begin
        saidaYMax<=123;
        saidaYm<=33;
    end
289:
    begin
        saidaYMax<=123;
        saidaYm<=33;
    end
290:
    begin
        saidaYMax<=123;
        saidaYm<=33;
    end
291:
    begin
        saidaYMax<=124;
        saidaYm<=34;
    end
292:
    begin
        saidaYMax<=124;
        saidaYm<=34;
    end
293:
    begin
        saidaYMax<=124;
        saidaYm<=34;
    end
294:
    begin
        saidaYMax<=124;
        saidaYm<=34;
    end
295:
    begin
        saidaYMax<=124;
        saidaYm<=34;
    end
296:
    begin
        saidaYMax<=124;
        saidaYm<=34;
    end
297:
    begin
        saidaYMax<=124;
        saidaYm<=34;
    end
298:
    begin
        saidaYMax<=124;
        saidaYm<=34;
    end
299:
    begin
        saidaYMax<=124;
        saidaYm<=34;
    end
300:
    begin
        saidaYMax<=124;
        saidaYm<=34;
    end
301:
    begin
        saidaYMax<=125;
        saidaYm<=35;
    end
302:
    begin
        saidaYMax<=125;
        saidaYm<=35;
    end
303:
    begin
        saidaYMax<=125;
        saidaYm<=35;
    end
304:
    begin
        saidaYMax<=125;
        saidaYm<=35;
    end
305:
    begin
        saidaYMax<=125;
        saidaYm<=35;
    end
306:
    begin
        saidaYMax<=125;
        saidaYm<=35;
    end
307:
    begin
        saidaYMax<=125;
        saidaYm<=35;
    end
308:
    begin
        saidaYMax<=125;
        saidaYm<=35;
    end
309:
    begin
        saidaYMax<=125;
        saidaYm<=35;
    end
310:
    begin
        saidaYMax<=125;
        saidaYm<=35;
    end
311:
    begin
        saidaYMax<=126;
        saidaYm<=36;
    end
312:
    begin
        saidaYMax<=126;
        saidaYm<=36;
    end
313:
    begin
        saidaYMax<=126;
        saidaYm<=36;
    end
314:
    begin
        saidaYMax<=126;
        saidaYm<=36;
    end
315:
    begin
        saidaYMax<=126;
        saidaYm<=36;
    end
316:
    begin
        saidaYMax<=126;
        saidaYm<=36;
    end
317:
    begin
        saidaYMax<=126;
        saidaYm<=36;
    end
318:
    begin
        saidaYMax<=126;
        saidaYm<=36;
    end
319:
    begin
        saidaYMax<=126;
        saidaYm<=36;
    end
320:
    begin
        saidaYMax<=126;
        saidaYm<=36;
    end
321:
    begin
        saidaYMax<=127;
        saidaYm<=37;
    end
322:
    begin
        saidaYMax<=127;
        saidaYm<=37;
    end
323:
    begin
        saidaYMax<=127;
        saidaYm<=37;
    end
324:
    begin
        saidaYMax<=127;
        saidaYm<=37;
    end
325:
    begin
        saidaYMax<=127;
        saidaYm<=37;
    end
326:
    begin
        saidaYMax<=127;
        saidaYm<=37;
    end
327:
    begin
        saidaYMax<=127;
        saidaYm<=37;
    end
328:
    begin
        saidaYMax<=127;
        saidaYm<=37;
    end
329:
    begin
        saidaYMax<=127;
        saidaYm<=37;
    end
330:
    begin
        saidaYMax<=127;
        saidaYm<=37;
    end
331:
    begin
        saidaYMax<=128;
        saidaYm<=38;
    end
332:
    begin
        saidaYMax<=128;
        saidaYm<=38;
    end
333:
    begin
        saidaYMax<=128;
        saidaYm<=38;
    end
334:
    begin
        saidaYMax<=128;
        saidaYm<=38;
    end
335:
    begin
        saidaYMax<=128;
        saidaYm<=38;
    end
336:
    begin
        saidaYMax<=128;
        saidaYm<=38;
    end
337:
    begin
        saidaYMax<=128;
        saidaYm<=38;
    end
338:
    begin
        saidaYMax<=128;
        saidaYm<=38;
    end
339:
    begin
        saidaYMax<=128;
        saidaYm<=38;
    end
340:
    begin
        saidaYMax<=128;
        saidaYm<=38;
    end
341:
    begin
        saidaYMax<=129;
        saidaYm<=39;
    end
342:
    begin
        saidaYMax<=129;
        saidaYm<=39;
    end
343:
    begin
        saidaYMax<=129;
        saidaYm<=39;
    end
344:
    begin
        saidaYMax<=129;
        saidaYm<=39;
    end
345:
    begin
        saidaYMax<=129;
        saidaYm<=39;
    end
346:
    begin
        saidaYMax<=129;
        saidaYm<=39;
    end
347:
    begin
        saidaYMax<=129;
        saidaYm<=39;
    end
348:
    begin
        saidaYMax<=129;
        saidaYm<=39;
    end
349:
    begin
        saidaYMax<=129;
        saidaYm<=39;
    end
350:
    begin
        saidaYMax<=129;
        saidaYm<=39;
    end
351:
    begin
        saidaYMax<=130;
        saidaYm<=40;
    end
352:
    begin
        saidaYMax<=130;
        saidaYm<=40;
    end
353:
    begin
        saidaYMax<=130;
        saidaYm<=40;
    end
354:
    begin
        saidaYMax<=130;
        saidaYm<=40;
    end
355:
    begin
        saidaYMax<=130;
        saidaYm<=40;
    end
356:
    begin
        saidaYMax<=130;
        saidaYm<=40;
    end
357:
    begin
        saidaYMax<=130;
        saidaYm<=40;
    end
358:
    begin
        saidaYMax<=130;
        saidaYm<=40;
    end
359:
    begin
        saidaYMax<=130;
        saidaYm<=40;
    end
360:
    begin
        saidaYMax<=130;
        saidaYm<=40;
    end
361:
    begin
        saidaYMax<=131;
        saidaYm<=41;
    end
362:
    begin
        saidaYMax<=131;
        saidaYm<=41;
    end
363:
    begin
        saidaYMax<=131;
        saidaYm<=41;
    end
364:
    begin
        saidaYMax<=131;
        saidaYm<=41;
    end
365:
    begin
        saidaYMax<=131;
        saidaYm<=41;
    end
366:
    begin
        saidaYMax<=131;
        saidaYm<=41;
    end
367:
    begin
        saidaYMax<=131;
        saidaYm<=41;
    end
368:
    begin
        saidaYMax<=131;
        saidaYm<=41;
    end
369:
    begin
        saidaYMax<=131;
        saidaYm<=41;
    end
370:
    begin
        saidaYMax<=131;
        saidaYm<=41;
    end
371:
    begin
        saidaYMax<=132;
        saidaYm<=42;
    end
372:
    begin
        saidaYMax<=132;
        saidaYm<=42;
    end
373:
    begin
        saidaYMax<=132;
        saidaYm<=42;
    end
374:
    begin
        saidaYMax<=132;
        saidaYm<=42;
    end
375:
    begin
        saidaYMax<=132;
        saidaYm<=42;
    end
376:
    begin
        saidaYMax<=132;
        saidaYm<=42;
    end
377:
    begin
        saidaYMax<=132;
        saidaYm<=42;
    end
378:
    begin
        saidaYMax<=132;
        saidaYm<=42;
    end
379:
    begin
        saidaYMax<=132;
        saidaYm<=42;
    end
380:
    begin
        saidaYMax<=132;
        saidaYm<=42;
    end
381:
    begin
        saidaYMax<=133;
        saidaYm<=43;
    end
382:
    begin
        saidaYMax<=133;
        saidaYm<=43;
    end
383:
    begin
        saidaYMax<=133;
        saidaYm<=43;
    end
384:
    begin
        saidaYMax<=133;
        saidaYm<=43;
    end
385:
    begin
        saidaYMax<=133;
        saidaYm<=43;
    end
386:
    begin
        saidaYMax<=133;
        saidaYm<=43;
    end
387:
    begin
        saidaYMax<=133;
        saidaYm<=43;
    end
388:
    begin
        saidaYMax<=133;
        saidaYm<=43;
    end
389:
    begin
        saidaYMax<=133;
        saidaYm<=43;
    end
390:
    begin
        saidaYMax<=133;
        saidaYm<=43;
    end
391:
    begin
        saidaYMax<=134;
        saidaYm<=44;
    end
392:
    begin
        saidaYMax<=134;
        saidaYm<=44;
    end
393:
    begin
        saidaYMax<=134;
        saidaYm<=44;
    end
394:
    begin
        saidaYMax<=134;
        saidaYm<=44;
    end
395:
    begin
        saidaYMax<=134;
        saidaYm<=44;
    end
396:
    begin
        saidaYMax<=134;
        saidaYm<=44;
    end
397:
    begin
        saidaYMax<=134;
        saidaYm<=44;
    end
398:
    begin
        saidaYMax<=134;
        saidaYm<=44;
    end
399:
    begin
        saidaYMax<=134;
        saidaYm<=44;
    end
400:
    begin
        saidaYMax<=134;
        saidaYm<=44;
    end
401:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
402:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
403:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
404:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
405:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
406:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
407:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
408:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
409:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
410:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
411:
    begin
        saidaYMax<=135;
        saidaYm<=45;
    end
412:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
413:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
414:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
415:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
416:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
417:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
418:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
419:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
420:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
421:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
422:
    begin
        saidaYMax<=136;
        saidaYm<=46;
    end
423:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
424:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
425:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
426:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
427:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
428:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
429:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
430:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
431:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
432:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
433:
    begin
        saidaYMax<=137;
        saidaYm<=47;
    end
434:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
435:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
436:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
437:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
438:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
439:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
440:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
441:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
442:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
443:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
444:
    begin
        saidaYMax<=138;
        saidaYm<=48;
    end
445:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
446:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
447:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
448:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
449:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
450:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
451:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
452:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
453:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
454:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
455:
    begin
        saidaYMax<=139;
        saidaYm<=49;
    end
456:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
457:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
458:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
459:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
460:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
461:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
462:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
463:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
464:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
465:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
466:
    begin
        saidaYMax<=140;
        saidaYm<=50;
    end
467:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
468:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
469:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
470:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
471:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
472:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
473:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
474:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
475:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
476:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
477:
    begin
        saidaYMax<=141;
        saidaYm<=51;
    end
478:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
479:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
480:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
481:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
482:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
483:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
484:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
485:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
486:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
487:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
488:
    begin
        saidaYMax<=142;
        saidaYm<=52;
    end
489:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
490:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
491:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
492:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
493:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
494:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
495:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
496:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
497:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
498:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
499:
    begin
        saidaYMax<=143;
        saidaYm<=53;
    end
500:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
501:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
502:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
503:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
504:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
505:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
506:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
507:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
508:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
509:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
510:
    begin
        saidaYMax<=144;
        saidaYm<=54;
    end
511:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
512:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
513:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
514:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
515:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
516:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
517:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
518:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
519:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
520:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
521:
    begin
        saidaYMax<=145;
        saidaYm<=55;
    end
522:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
523:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
524:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
525:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
526:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
527:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
528:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
529:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
530:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
531:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
532:
    begin
        saidaYMax<=146;
        saidaYm<=56;
    end
533:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
534:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
535:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
536:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
537:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
538:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
539:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
540:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
541:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
542:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
543:
    begin
        saidaYMax<=147;
        saidaYm<=57;
    end
544:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
545:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
546:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
547:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
548:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
549:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
550:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
551:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
552:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
553:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
554:
    begin
        saidaYMax<=148;
        saidaYm<=58;
    end
555:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
556:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
557:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
558:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
559:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
560:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
561:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
562:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
563:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
564:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
565:
    begin
        saidaYMax<=149;
        saidaYm<=59;
    end
566:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
567:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
568:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
569:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
570:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
571:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
572:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
573:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
574:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
575:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
576:
    begin
        saidaYMax<=150;
        saidaYm<=60;
    end
577:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
578:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
579:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
580:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
581:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
582:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
583:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
584:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
585:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
586:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
587:
    begin
        saidaYMax<=151;
        saidaYm<=61;
    end
588:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
589:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
590:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
591:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
592:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
593:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
594:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
595:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
596:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
597:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
598:
    begin
        saidaYMax<=152;
        saidaYm<=62;
    end
599:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
600:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
601:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
602:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
603:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
604:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
605:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
606:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
607:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
608:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
609:
    begin
        saidaYMax<=153;
        saidaYm<=63;
    end
610:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
611:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
612:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
613:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
614:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
615:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
616:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
617:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
618:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
619:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
620:
    begin
        saidaYMax<=154;
        saidaYm<=64;
    end
621:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
622:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
623:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
624:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
625:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
626:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
627:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
628:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
629:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
630:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
631:
    begin
        saidaYMax<=155;
        saidaYm<=65;
    end
632:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
633:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
634:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
635:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
636:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
637:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
638:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
639:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
640:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
641:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
642:
    begin
        saidaYMax<=156;
        saidaYm<=66;
    end
643:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
644:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
645:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
646:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
647:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
648:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
649:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
650:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
651:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
652:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
653:
    begin
        saidaYMax<=157;
        saidaYm<=67;
    end
654:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
655:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
656:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
657:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
658:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
659:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
660:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
661:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
662:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
663:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
664:
    begin
        saidaYMax<=158;
        saidaYm<=68;
    end
665:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
666:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
667:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
668:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
669:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
670:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
671:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
672:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
673:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
674:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
675:
    begin
        saidaYMax<=159;
        saidaYm<=69;
    end
676:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
677:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
678:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
679:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
680:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
681:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
682:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
683:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
684:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
685:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
686:
    begin
        saidaYMax<=160;
        saidaYm<=70;
    end
687:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
688:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
689:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
690:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
691:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
692:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
693:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
694:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
695:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
696:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
697:
    begin
        saidaYMax<=161;
        saidaYm<=71;
    end
698:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
699:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
700:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
701:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
702:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
703:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
704:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
705:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
706:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
707:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
708:
    begin
        saidaYMax<=162;
        saidaYm<=72;
    end
709:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
710:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
711:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
712:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
713:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
714:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
715:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
716:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
717:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
718:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
719:
    begin
        saidaYMax<=163;
        saidaYm<=73;
    end
720:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
721:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
722:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
723:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
724:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
725:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
726:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
727:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
728:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
729:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
730:
    begin
        saidaYMax<=164;
        saidaYm<=74;
    end
731:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
732:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
733:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
734:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
735:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
736:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
737:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
738:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
739:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
740:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
741:
    begin
        saidaYMax<=165;
        saidaYm<=75;
    end
742:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
743:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
744:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
745:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
746:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
747:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
748:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
749:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
750:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
751:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
752:
    begin
        saidaYMax<=166;
        saidaYm<=76;
    end
753:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
754:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
755:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
756:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
757:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
758:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
759:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
760:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
761:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
762:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
763:
    begin
        saidaYMax<=167;
        saidaYm<=77;
    end
764:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
765:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
766:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
767:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
768:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
769:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
770:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
771:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
772:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
773:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
774:
    begin
        saidaYMax<=168;
        saidaYm<=78;
    end
775:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
776:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
777:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
778:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
779:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
780:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
781:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
782:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
783:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
784:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
785:
    begin
        saidaYMax<=169;
        saidaYm<=79;
    end
786:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
787:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
788:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
789:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
790:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
791:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
792:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
793:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
794:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
795:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
796:
    begin
        saidaYMax<=170;
        saidaYm<=80;
    end
797:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
798:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
799:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
800:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
801:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
802:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
803:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
804:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
805:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
806:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
807:
    begin
        saidaYMax<=171;
        saidaYm<=81;
    end
808:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
809:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
810:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
811:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
812:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
813:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
814:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
815:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
816:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
817:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
818:
    begin
        saidaYMax<=172;
        saidaYm<=82;
    end
819:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
820:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
821:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
822:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
823:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
824:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
825:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
826:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
827:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
828:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
829:
    begin
        saidaYMax<=173;
        saidaYm<=83;
    end
830:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
831:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
832:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
833:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
834:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
835:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
836:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
837:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
838:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
839:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
840:
    begin
        saidaYMax<=174;
        saidaYm<=84;
    end
841:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
842:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
843:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
844:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
845:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
846:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
847:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
848:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
849:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
850:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
851:
    begin
        saidaYMax<=175;
        saidaYm<=85;
    end
852:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
853:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
854:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
855:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
856:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
857:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
858:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
859:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
860:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
861:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
862:
    begin
        saidaYMax<=176;
        saidaYm<=86;
    end
863:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
864:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
865:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
866:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
867:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
868:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
869:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
870:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
871:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
872:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
873:
    begin
        saidaYMax<=177;
        saidaYm<=87;
    end
874:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
875:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
876:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
877:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
878:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
879:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
880:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
881:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
882:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
883:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
884:
    begin
        saidaYMax<=178;
        saidaYm<=88;
    end
885:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
886:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
887:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
888:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
889:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
890:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
891:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
892:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
893:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
894:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
895:
    begin
        saidaYMax<=179;
        saidaYm<=89;
    end
896:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
897:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
898:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
899:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
900:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
901:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
902:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
903:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
904:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
905:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
906:
    begin
        saidaYMax<=180;
        saidaYm<=90;
    end
907:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
908:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
909:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
910:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
911:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
912:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
913:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
914:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
915:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
916:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
917:
    begin
        saidaYMax<=181;
        saidaYm<=91;
    end
918:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
919:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
920:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
921:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
922:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
923:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
924:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
925:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
926:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
927:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
928:
    begin
        saidaYMax<=182;
        saidaYm<=92;
    end
929:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
930:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
931:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
932:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
933:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
934:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
935:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
936:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
937:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
938:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
939:
    begin
        saidaYMax<=183;
        saidaYm<=93;
    end
940:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
941:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
942:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
943:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
944:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
945:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
946:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
947:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
948:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
949:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
950:
    begin
        saidaYMax<=184;
        saidaYm<=94;
    end
951:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
952:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
953:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
954:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
955:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
956:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
957:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
958:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
959:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
960:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
961:
    begin
        saidaYMax<=185;
        saidaYm<=95;
    end
962:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
963:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
964:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
965:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
966:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
967:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
968:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
969:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
970:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
971:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
972:
    begin
        saidaYMax<=186;
        saidaYm<=96;
    end
973:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
974:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
975:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
976:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
977:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
978:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
979:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
980:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
981:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
982:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
983:
    begin
        saidaYMax<=187;
        saidaYm<=97;
    end
984:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
985:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
986:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
987:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
988:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
989:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
990:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
991:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
992:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
993:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
994:
    begin
        saidaYMax<=188;
        saidaYm<=98;
    end
995:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
996:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
997:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
998:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
999:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
1000:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
1001:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
1002:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
1003:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
1004:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
1005:
    begin
        saidaYMax<=189;
        saidaYm<=99;
    end
1006:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1007:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1008:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1009:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1010:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1011:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1012:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1013:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1014:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1015:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1016:
    begin
        saidaYMax<=190;
        saidaYm<=100;
    end
1017:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1018:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1019:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1020:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1021:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1022:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1023:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1024:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1025:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1026:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1027:
    begin
        saidaYMax<=191;
        saidaYm<=101;
    end
1028:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1029:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1030:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1031:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1032:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1033:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1034:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1035:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1036:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1037:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1038:
    begin
        saidaYMax<=192;
        saidaYm<=102;
    end
1039:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1040:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1041:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1042:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1043:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1044:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1045:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1046:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1047:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1048:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1049:
    begin
        saidaYMax<=193;
        saidaYm<=103;
    end
1050:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1051:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1052:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1053:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1054:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1055:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1056:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1057:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1058:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1059:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1060:
    begin
        saidaYMax<=194;
        saidaYm<=104;
    end
1061:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1062:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1063:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1064:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1065:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1066:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1067:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1068:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1069:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1070:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1071:
    begin
        saidaYMax<=195;
        saidaYm<=105;
    end
1072:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1073:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1074:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1075:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1076:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1077:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1078:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1079:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1080:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1081:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1082:
    begin
        saidaYMax<=196;
        saidaYm<=106;
    end
1083:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1084:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1085:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1086:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1087:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1088:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1089:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1090:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1091:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1092:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1093:
    begin
        saidaYMax<=197;
        saidaYm<=107;
    end
1094:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1095:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1096:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1097:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1098:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1099:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1100:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1101:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1102:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1103:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1104:
    begin
        saidaYMax<=198;
        saidaYm<=108;
    end
1105:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1106:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1107:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1108:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1109:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1110:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1111:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1112:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1113:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1114:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1115:
    begin
        saidaYMax<=199;
        saidaYm<=109;
    end
1116:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1117:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1118:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1119:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1120:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1121:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1122:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1123:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1124:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1125:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1126:
    begin
        saidaYMax<=200;
        saidaYm<=110;
    end
1127:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1128:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1129:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1130:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1131:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1132:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1133:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1134:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1135:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1136:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1137:
    begin
        saidaYMax<=201;
        saidaYm<=111;
    end
1138:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1139:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1140:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1141:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1142:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1143:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1144:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1145:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1146:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1147:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1148:
    begin
        saidaYMax<=202;
        saidaYm<=112;
    end
1149:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1150:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1151:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1152:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1153:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1154:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1155:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1156:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1157:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1158:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1159:
    begin
        saidaYMax<=203;
        saidaYm<=113;
    end
1160:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1161:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1162:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1163:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1164:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1165:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1166:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1167:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1168:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1169:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1170:
    begin
        saidaYMax<=204;
        saidaYm<=114;
    end
1171:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1172:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1173:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1174:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1175:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1176:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1177:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1178:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1179:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1180:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1181:
    begin
        saidaYMax<=205;
        saidaYm<=115;
    end
1182:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1183:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1184:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1185:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1186:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1187:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1188:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1189:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1190:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1191:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1192:
    begin
        saidaYMax<=206;
        saidaYm<=116;
    end
1193:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1194:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1195:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1196:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1197:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1198:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1199:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1200:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1201:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1202:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1203:
    begin
        saidaYMax<=207;
        saidaYm<=117;
    end
1204:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1205:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1206:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1207:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1208:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1209:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1210:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1211:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1212:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1213:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1214:
    begin
        saidaYMax<=208;
        saidaYm<=118;
    end
1215:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1216:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1217:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1218:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1219:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1220:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1221:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1222:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1223:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1224:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1225:
    begin
        saidaYMax<=209;
        saidaYm<=119;
    end
1226:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1227:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1228:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1229:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1230:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1231:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1232:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1233:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1234:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1235:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1236:
    begin
        saidaYMax<=210;
        saidaYm<=120;
    end
1237:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1238:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1239:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1240:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1241:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1242:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1243:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1244:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1245:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1246:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1247:
    begin
        saidaYMax<=211;
        saidaYm<=121;
    end
1248:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1249:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1250:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1251:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1252:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1253:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1254:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1255:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1256:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1257:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1258:
    begin
        saidaYMax<=212;
        saidaYm<=122;
    end
1259:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1260:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1261:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1262:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1263:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1264:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1265:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1266:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1267:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1268:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1269:
    begin
        saidaYMax<=213;
        saidaYm<=123;
    end
1270:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1271:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1272:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1273:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1274:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1275:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1276:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1277:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1278:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1279:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1280:
    begin
        saidaYMax<=214;
        saidaYm<=124;
    end
1281:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1282:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1283:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1284:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1285:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1286:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1287:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1288:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1289:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1290:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1291:
    begin
        saidaYMax<=215;
        saidaYm<=125;
    end
1292:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1293:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1294:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1295:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1296:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1297:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1298:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1299:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1300:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1301:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1302:
    begin
        saidaYMax<=216;
        saidaYm<=126;
    end
1303:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1304:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1305:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1306:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1307:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1308:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1309:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1310:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1311:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1312:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1313:
    begin
        saidaYMax<=217;
        saidaYm<=127;
    end
1314:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1315:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1316:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1317:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1318:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1319:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1320:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1321:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1322:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1323:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1324:
    begin
        saidaYMax<=218;
        saidaYm<=128;
    end
1325:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1326:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1327:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1328:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1329:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1330:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1331:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1332:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1333:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1334:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1335:
    begin
        saidaYMax<=219;
        saidaYm<=129;
    end
1336:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1337:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1338:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1339:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1340:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1341:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1342:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1343:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1344:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1345:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1346:
    begin
        saidaYMax<=220;
        saidaYm<=130;
    end
1347:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1348:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1349:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1350:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1351:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1352:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1353:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1354:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1355:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1356:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1357:
    begin
        saidaYMax<=221;
        saidaYm<=131;
    end
1358:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1359:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1360:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1361:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1362:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1363:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1364:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1365:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1366:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1367:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1368:
    begin
        saidaYMax<=222;
        saidaYm<=132;
    end
1369:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1370:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1371:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1372:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1373:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1374:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1375:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1376:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1377:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1378:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1379:
    begin
        saidaYMax<=223;
        saidaYm<=133;
    end
1380:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1381:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1382:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1383:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1384:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1385:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1386:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1387:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1388:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1389:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1390:
    begin
        saidaYMax<=224;
        saidaYm<=134;
    end
1391:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1392:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1393:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1394:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1395:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1396:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1397:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1398:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1399:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1400:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1401:
    begin
        saidaYMax<=225;
        saidaYm<=135;
    end
1402:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1403:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1404:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1405:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1406:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1407:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1408:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1409:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1410:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1411:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1412:
    begin
        saidaYMax<=226;
        saidaYm<=136;
    end
1413:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1414:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1415:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1416:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1417:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1418:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1419:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1420:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1421:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1422:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1423:
    begin
        saidaYMax<=227;
        saidaYm<=137;
    end
1424:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1425:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1426:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1427:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1428:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1429:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1430:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1431:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1432:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1433:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1434:
    begin
        saidaYMax<=228;
        saidaYm<=138;
    end
1435:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1436:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1437:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1438:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1439:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1440:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1441:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1442:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1443:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1444:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1445:
    begin
        saidaYMax<=229;
        saidaYm<=139;
    end
1446:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1447:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1448:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1449:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1450:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1451:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1452:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1453:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1454:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1455:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1456:
    begin
        saidaYMax<=230;
        saidaYm<=140;
    end
1457:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1458:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1459:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1460:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1461:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1462:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1463:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1464:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1465:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1466:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1467:
    begin
        saidaYMax<=231;
        saidaYm<=141;
    end
1468:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1469:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1470:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1471:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1472:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1473:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1474:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1475:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1476:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1477:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1478:
    begin
        saidaYMax<=232;
        saidaYm<=142;
    end
1479:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1480:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1481:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1482:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1483:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1484:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1485:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1486:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1487:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1488:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1489:
    begin
        saidaYMax<=233;
        saidaYm<=143;
    end
1490:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1491:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1492:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1493:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1494:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1495:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1496:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1497:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1498:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1499:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1500:
    begin
        saidaYMax<=234;
        saidaYm<=144;
    end
1501:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1502:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1503:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1504:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1505:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1506:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1507:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1508:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1509:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1510:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1511:
    begin
        saidaYMax<=235;
        saidaYm<=145;
    end
1512:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1513:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1514:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1515:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1516:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1517:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1518:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1519:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1520:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1521:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1522:
    begin
        saidaYMax<=236;
        saidaYm<=146;
    end
1523:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1524:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1525:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1526:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1527:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1528:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1529:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1530:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1531:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1532:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1533:
    begin
        saidaYMax<=237;
        saidaYm<=147;
    end
1534:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1535:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1536:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1537:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1538:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1539:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1540:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1541:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1542:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1543:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1544:
    begin
        saidaYMax<=238;
        saidaYm<=148;
    end
1545:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1546:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1547:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1548:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1549:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1550:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1551:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1552:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1553:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1554:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1555:
    begin
        saidaYMax<=239;
        saidaYm<=149;
    end
1556:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1557:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1558:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1559:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1560:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1561:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1562:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1563:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1564:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1565:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1566:
    begin
        saidaYMax<=240;
        saidaYm<=150;
    end
1567:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1568:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1569:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1570:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1571:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1572:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1573:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1574:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1575:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1576:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1577:
    begin
        saidaYMax<=241;
        saidaYm<=151;
    end
1578:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1579:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1580:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1581:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1582:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1583:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1584:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1585:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1586:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1587:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1588:
    begin
        saidaYMax<=242;
        saidaYm<=152;
    end
1589:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1590:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1591:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1592:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1593:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1594:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1595:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1596:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1597:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1598:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1599:
    begin
        saidaYMax<=243;
        saidaYm<=153;
    end
1600:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1601:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1602:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1603:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1604:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1605:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1606:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1607:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1608:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1609:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1610:
    begin
        saidaYMax<=244;
        saidaYm<=154;
    end
1611:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1612:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1613:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1614:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1615:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1616:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1617:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1618:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1619:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1620:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1621:
    begin
        saidaYMax<=245;
        saidaYm<=155;
    end
1622:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1623:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1624:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1625:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1626:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1627:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1628:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1629:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1630:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1631:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1632:
    begin
        saidaYMax<=246;
        saidaYm<=156;
    end
1633:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1634:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1635:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1636:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1637:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1638:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1639:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1640:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1641:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1642:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1643:
    begin
        saidaYMax<=247;
        saidaYm<=157;
    end
1644:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1645:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1646:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1647:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1648:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1649:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1650:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1651:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1652:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1653:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1654:
    begin
        saidaYMax<=248;
        saidaYm<=158;
    end
1655:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1656:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1657:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1658:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1659:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1660:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1661:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1662:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1663:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1664:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1665:
    begin
        saidaYMax<=249;
        saidaYm<=159;
    end
1666:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1667:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1668:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1669:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1670:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1671:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1672:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1673:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1674:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1675:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1676:
    begin
        saidaYMax<=250;
        saidaYm<=160;
    end
1677:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1678:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1679:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1680:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1681:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1682:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1683:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1684:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1685:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1686:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1687:
    begin
        saidaYMax<=251;
        saidaYm<=161;
    end
1688:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1689:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1690:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1691:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1692:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1693:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1694:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1695:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1696:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1697:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1698:
    begin
        saidaYMax<=252;
        saidaYm<=162;
    end
1699:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1700:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1701:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1702:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1703:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1704:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1705:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1706:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1707:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1708:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1709:
    begin
        saidaYMax<=253;
        saidaYm<=163;
    end
1710:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1711:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1712:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1713:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1714:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1715:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1716:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1717:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1718:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1719:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1720:
    begin
        saidaYMax<=254;
        saidaYm<=164;
    end
1721:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1722:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1723:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1724:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1725:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1726:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1727:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1728:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1729:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1730:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1731:
    begin
        saidaYMax<=255;
        saidaYm<=165;
    end
1732:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1733:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1734:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1735:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1736:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1737:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1738:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1739:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1740:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1741:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1742:
    begin
        saidaYMax<=256;
        saidaYm<=166;
    end
1743:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1744:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1745:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1746:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1747:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1748:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1749:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1750:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1751:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1752:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1753:
    begin
        saidaYMax<=257;
        saidaYm<=167;
    end
1754:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1755:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1756:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1757:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1758:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1759:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1760:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1761:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1762:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1763:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1764:
    begin
        saidaYMax<=258;
        saidaYm<=168;
    end
1765:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1766:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1767:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1768:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1769:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1770:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1771:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1772:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1773:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1774:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1775:
    begin
        saidaYMax<=259;
        saidaYm<=169;
    end
1776:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1777:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1778:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1779:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1780:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1781:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1782:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1783:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1784:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1785:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1786:
    begin
        saidaYMax<=260;
        saidaYm<=170;
    end
1787:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1788:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1789:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1790:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1791:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1792:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1793:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1794:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1795:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1796:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1797:
    begin
        saidaYMax<=261;
        saidaYm<=171;
    end
1798:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1799:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1800:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1801:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1802:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1803:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1804:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1805:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1806:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1807:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1808:
    begin
        saidaYMax<=262;
        saidaYm<=172;
    end
1809:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1810:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1811:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1812:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1813:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1814:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1815:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1816:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1817:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1818:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1819:
    begin
        saidaYMax<=263;
        saidaYm<=173;
    end
1820:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1821:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1822:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1823:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1824:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1825:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1826:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1827:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1828:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1829:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1830:
    begin
        saidaYMax<=264;
        saidaYm<=174;
    end
1831:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1832:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1833:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1834:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1835:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1836:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1837:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1838:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1839:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1840:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1841:
    begin
        saidaYMax<=265;
        saidaYm<=175;
    end
1842:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1843:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1844:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1845:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1846:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1847:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1848:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1849:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1850:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1851:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1852:
    begin
        saidaYMax<=266;
        saidaYm<=176;
    end
1853:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1854:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1855:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1856:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1857:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1858:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1859:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1860:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1861:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1862:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1863:
    begin
        saidaYMax<=267;
        saidaYm<=177;
    end
1864:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1865:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1866:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1867:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1868:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1869:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1870:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1871:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1872:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1873:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1874:
    begin
        saidaYMax<=268;
        saidaYm<=178;
    end
1875:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1876:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1877:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1878:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1879:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1880:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1881:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1882:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1883:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1884:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1885:
    begin
        saidaYMax<=269;
        saidaYm<=179;
    end
1886:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1887:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1888:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1889:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1890:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1891:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1892:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1893:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1894:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1895:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1896:
    begin
        saidaYMax<=270;
        saidaYm<=180;
    end
1897:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1898:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1899:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1900:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1901:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1902:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1903:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1904:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1905:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1906:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1907:
    begin
        saidaYMax<=271;
        saidaYm<=181;
    end
1908:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1909:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1910:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1911:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1912:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1913:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1914:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1915:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1916:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1917:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1918:
    begin
        saidaYMax<=272;
        saidaYm<=182;
    end
1919:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1920:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1921:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1922:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1923:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1924:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1925:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1926:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1927:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1928:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1929:
    begin
        saidaYMax<=273;
        saidaYm<=183;
    end
1930:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1931:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1932:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1933:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1934:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1935:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1936:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1937:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1938:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1939:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1940:
    begin
        saidaYMax<=274;
        saidaYm<=184;
    end
1941:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1942:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1943:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1944:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1945:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1946:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1947:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1948:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1949:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1950:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1951:
    begin
        saidaYMax<=275;
        saidaYm<=185;
    end
1952:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1953:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1954:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1955:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1956:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1957:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1958:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1959:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1960:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1961:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1962:
    begin
        saidaYMax<=276;
        saidaYm<=186;
    end
1963:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1964:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1965:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1966:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1967:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1968:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1969:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1970:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1971:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1972:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1973:
    begin
        saidaYMax<=277;
        saidaYm<=187;
    end
1974:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1975:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1976:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1977:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1978:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1979:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1980:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1981:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1982:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1983:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1984:
    begin
        saidaYMax<=278;
        saidaYm<=188;
    end
1985:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1986:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1987:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1988:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1989:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1990:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1991:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1992:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1993:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1994:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1995:
    begin
        saidaYMax<=279;
        saidaYm<=189;
    end
1996:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
1997:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
1998:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
1999:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
2000:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
2001:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
2002:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
2003:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
2004:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
2005:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
2006:
    begin
        saidaYMax<=280;
        saidaYm<=190;
    end
2007:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2008:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2009:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2010:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2011:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2012:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2013:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2014:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2015:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2016:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2017:
    begin
        saidaYMax<=281;
        saidaYm<=191;
    end
2018:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2019:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2020:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2021:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2022:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2023:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2024:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2025:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2026:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2027:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2028:
    begin
        saidaYMax<=282;
        saidaYm<=192;
    end
2029:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2030:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2031:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2032:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2033:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2034:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2035:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2036:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2037:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2038:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2039:
    begin
        saidaYMax<=283;
        saidaYm<=193;
    end
2040:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2041:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2042:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2043:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2044:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2045:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2046:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2047:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2048:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2049:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2050:
    begin
        saidaYMax<=284;
        saidaYm<=194;
    end
2051:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2052:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2053:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2054:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2055:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2056:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2057:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2058:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2059:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2060:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2061:
    begin
        saidaYMax<=285;
        saidaYm<=195;
    end
2062:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2063:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2064:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2065:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2066:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2067:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2068:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2069:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2070:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2071:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2072:
    begin
        saidaYMax<=286;
        saidaYm<=196;
    end
2073:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2074:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2075:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2076:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2077:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2078:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2079:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2080:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2081:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2082:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2083:
    begin
        saidaYMax<=287;
        saidaYm<=197;
    end
2084:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2085:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2086:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2087:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2088:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2089:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2090:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2091:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2092:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2093:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2094:
    begin
        saidaYMax<=288;
        saidaYm<=198;
    end
2095:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2096:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2097:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2098:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2099:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2100:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2101:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2102:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2103:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2104:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2105:
    begin
        saidaYMax<=289;
        saidaYm<=199;
    end
2106:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2107:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2108:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2109:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2110:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2111:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2112:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2113:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2114:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2115:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2116:
    begin
        saidaYMax<=290;
        saidaYm<=200;
    end
2117:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2118:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2119:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2120:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2121:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2122:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2123:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2124:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2125:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2126:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2127:
    begin
        saidaYMax<=291;
        saidaYm<=201;
    end
2128:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2129:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2130:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2131:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2132:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2133:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2134:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2135:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2136:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2137:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2138:
    begin
        saidaYMax<=292;
        saidaYm<=202;
    end
2139:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2140:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2141:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2142:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2143:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2144:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2145:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2146:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2147:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2148:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2149:
    begin
        saidaYMax<=293;
        saidaYm<=203;
    end
2150:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2151:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2152:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2153:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2154:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2155:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2156:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2157:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2158:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2159:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2160:
    begin
        saidaYMax<=294;
        saidaYm<=204;
    end
2161:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2162:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2163:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2164:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2165:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2166:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2167:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2168:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2169:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2170:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2171:
    begin
        saidaYMax<=295;
        saidaYm<=205;
    end
2172:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2173:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2174:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2175:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2176:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2177:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2178:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2179:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2180:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2181:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2182:
    begin
        saidaYMax<=296;
        saidaYm<=206;
    end
2183:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2184:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2185:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2186:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2187:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2188:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2189:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2190:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2191:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2192:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2193:
    begin
        saidaYMax<=297;
        saidaYm<=207;
    end
2194:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2195:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2196:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2197:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2198:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2199:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2200:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2201:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2202:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2203:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2204:
    begin
        saidaYMax<=298;
        saidaYm<=208;
    end
2205:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2206:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2207:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2208:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2209:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2210:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2211:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2212:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2213:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2214:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2215:
    begin
        saidaYMax<=299;
        saidaYm<=209;
    end
2216:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2217:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2218:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2219:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2220:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2221:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2222:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2223:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2224:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2225:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2226:
    begin
        saidaYMax<=300;
        saidaYm<=210;
    end
2227:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2228:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2229:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2230:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2231:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2232:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2233:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2234:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2235:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2236:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2237:
    begin
        saidaYMax<=301;
        saidaYm<=211;
    end
2238:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2239:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2240:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2241:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2242:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2243:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2244:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2245:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2246:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2247:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2248:
    begin
        saidaYMax<=302;
        saidaYm<=212;
    end
2249:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2250:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2251:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2252:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2253:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2254:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2255:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2256:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2257:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2258:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2259:
    begin
        saidaYMax<=303;
        saidaYm<=213;
    end
2260:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2261:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2262:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2263:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2264:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2265:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2266:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2267:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2268:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2269:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2270:
    begin
        saidaYMax<=304;
        saidaYm<=214;
    end
2271:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2272:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2273:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2274:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2275:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2276:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2277:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2278:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2279:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2280:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2281:
    begin
        saidaYMax<=305;
        saidaYm<=215;
    end
2282:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2283:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2284:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2285:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2286:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2287:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2288:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2289:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2290:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2291:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2292:
    begin
        saidaYMax<=306;
        saidaYm<=216;
    end
2293:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2294:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2295:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2296:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2297:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2298:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2299:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2300:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2301:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2302:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2303:
    begin
        saidaYMax<=307;
        saidaYm<=217;
    end
2304:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2305:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2306:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2307:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2308:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2309:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2310:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2311:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2312:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2313:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2314:
    begin
        saidaYMax<=308;
        saidaYm<=218;
    end
2315:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2316:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2317:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2318:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2319:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2320:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2321:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2322:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2323:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2324:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2325:
    begin
        saidaYMax<=309;
        saidaYm<=219;
    end
2326:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2327:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2328:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2329:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2330:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2331:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2332:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2333:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2334:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2335:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2336:
    begin
        saidaYMax<=310;
        saidaYm<=220;
    end
2337:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2338:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2339:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2340:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2341:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2342:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2343:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2344:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2345:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2346:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2347:
    begin
        saidaYMax<=311;
        saidaYm<=221;
    end
2348:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2349:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2350:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2351:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2352:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2353:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2354:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2355:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2356:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2357:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2358:
    begin
        saidaYMax<=312;
        saidaYm<=222;
    end
2359:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2360:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2361:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2362:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2363:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2364:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2365:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2366:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2367:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2368:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2369:
    begin
        saidaYMax<=313;
        saidaYm<=223;
    end
2370:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2371:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2372:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2373:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2374:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2375:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2376:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2377:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2378:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2379:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2380:
    begin
        saidaYMax<=314;
        saidaYm<=224;
    end
2381:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2382:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2383:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2384:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2385:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2386:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2387:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2388:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2389:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2390:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2391:
    begin
        saidaYMax<=315;
        saidaYm<=225;
    end
2392:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2393:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2394:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2395:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2396:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2397:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2398:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2399:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2400:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2401:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2402:
    begin
        saidaYMax<=316;
        saidaYm<=226;
    end
2403:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2404:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2405:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2406:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2407:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2408:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2409:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2410:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2411:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2412:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2413:
    begin
        saidaYMax<=317;
        saidaYm<=227;
    end
2414:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2415:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2416:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2417:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2418:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2419:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2420:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2421:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2422:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2423:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2424:
    begin
        saidaYMax<=318;
        saidaYm<=228;
    end
2425:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2426:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2427:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2428:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2429:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2430:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2431:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2432:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2433:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2434:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2435:
    begin
        saidaYMax<=319;
        saidaYm<=229;
    end
2436:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2437:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2438:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2439:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2440:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2441:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2442:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2443:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2444:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2445:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2446:
    begin
        saidaYMax<=320;
        saidaYm<=230;
    end
2447:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2448:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2449:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2450:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2451:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2452:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2453:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2454:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2455:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2456:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2457:
    begin
        saidaYMax<=321;
        saidaYm<=231;
    end
2458:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2459:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2460:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2461:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2462:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2463:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2464:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2465:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2466:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2467:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2468:
    begin
        saidaYMax<=322;
        saidaYm<=232;
    end
2469:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2470:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2471:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2472:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2473:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2474:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2475:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2476:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2477:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2478:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2479:
    begin
        saidaYMax<=323;
        saidaYm<=233;
    end
2480:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2481:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2482:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2483:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2484:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2485:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2486:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2487:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2488:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2489:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2490:
    begin
        saidaYMax<=324;
        saidaYm<=234;
    end
2491:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2492:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2493:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2494:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2495:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2496:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2497:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2498:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2499:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2500:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2501:
    begin
        saidaYMax<=325;
        saidaYm<=235;
    end
2502:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2503:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2504:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2505:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2506:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2507:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2508:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2509:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2510:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2511:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2512:
    begin
        saidaYMax<=326;
        saidaYm<=236;
    end
2513:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2514:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2515:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2516:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2517:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2518:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2519:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2520:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2521:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2522:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2523:
    begin
        saidaYMax<=327;
        saidaYm<=237;
    end
2524:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2525:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2526:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2527:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2528:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2529:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2530:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2531:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2532:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2533:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2534:
    begin
        saidaYMax<=328;
        saidaYm<=238;
    end
2535:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2536:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2537:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2538:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2539:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2540:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2541:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2542:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2543:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2544:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2545:
    begin
        saidaYMax<=329;
        saidaYm<=239;
    end
2546:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2547:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2548:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2549:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2550:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2551:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2552:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2553:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2554:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2555:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2556:
    begin
        saidaYMax<=330;
        saidaYm<=240;
    end
2557:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2558:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2559:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2560:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2561:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2562:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2563:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2564:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2565:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2566:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2567:
    begin
        saidaYMax<=331;
        saidaYm<=241;
    end
2568:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2569:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2570:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2571:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2572:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2573:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2574:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2575:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2576:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2577:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2578:
    begin
        saidaYMax<=332;
        saidaYm<=242;
    end
2579:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2580:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2581:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2582:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2583:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2584:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2585:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2586:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2587:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2588:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2589:
    begin
        saidaYMax<=333;
        saidaYm<=243;
    end
2590:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2591:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2592:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2593:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2594:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2595:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2596:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2597:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2598:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2599:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2600:
    begin
        saidaYMax<=334;
        saidaYm<=244;
    end
2601:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2602:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2603:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2604:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2605:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2606:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2607:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2608:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2609:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2610:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2611:
    begin
        saidaYMax<=335;
        saidaYm<=245;
    end
2612:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2613:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2614:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2615:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2616:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2617:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2618:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2619:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2620:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2621:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2622:
    begin
        saidaYMax<=336;
        saidaYm<=246;
    end
2623:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2624:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2625:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2626:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2627:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2628:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2629:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2630:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2631:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2632:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2633:
    begin
        saidaYMax<=337;
        saidaYm<=247;
    end
2634:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2635:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2636:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2637:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2638:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2639:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2640:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2641:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2642:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2643:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2644:
    begin
        saidaYMax<=338;
        saidaYm<=248;
    end
2645:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2646:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2647:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2648:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2649:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2650:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2651:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2652:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2653:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2654:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2655:
    begin
        saidaYMax<=339;
        saidaYm<=249;
    end
2656:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2657:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2658:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2659:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2660:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2661:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2662:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2663:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2664:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2665:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2666:
    begin
        saidaYMax<=340;
        saidaYm<=250;
    end
2667:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2668:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2669:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2670:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2671:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2672:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2673:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2674:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2675:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2676:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2677:
    begin
        saidaYMax<=341;
        saidaYm<=251;
    end
2678:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2679:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2680:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2681:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2682:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2683:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2684:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2685:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2686:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2687:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2688:
    begin
        saidaYMax<=342;
        saidaYm<=252;
    end
2689:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2690:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2691:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2692:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2693:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2694:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2695:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2696:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2697:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2698:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2699:
    begin
        saidaYMax<=343;
        saidaYm<=253;
    end
2700:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2701:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2702:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2703:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2704:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2705:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2706:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2707:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2708:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2709:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2710:
    begin
        saidaYMax<=344;
        saidaYm<=254;
    end
2711:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2712:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2713:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2714:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2715:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2716:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2717:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2718:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2719:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2720:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2721:
    begin
        saidaYMax<=345;
        saidaYm<=255;
    end
2722:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2723:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2724:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2725:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2726:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2727:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2728:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2729:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2730:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2731:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2732:
    begin
        saidaYMax<=346;
        saidaYm<=256;
    end
2733:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2734:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2735:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2736:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2737:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2738:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2739:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2740:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2741:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2742:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2743:
    begin
        saidaYMax<=347;
        saidaYm<=257;
    end
2744:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2745:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2746:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2747:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2748:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2749:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2750:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2751:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2752:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2753:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2754:
    begin
        saidaYMax<=348;
        saidaYm<=258;
    end
2755:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2756:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2757:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2758:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2759:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2760:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2761:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2762:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2763:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2764:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2765:
    begin
        saidaYMax<=349;
        saidaYm<=259;
    end
2766:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2767:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2768:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2769:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2770:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2771:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2772:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2773:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2774:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2775:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2776:
    begin
        saidaYMax<=350;
        saidaYm<=260;
    end
2777:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2778:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2779:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2780:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2781:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2782:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2783:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2784:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2785:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2786:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2787:
    begin
        saidaYMax<=351;
        saidaYm<=261;
    end
2788:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2789:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2790:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2791:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2792:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2793:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2794:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2795:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2796:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2797:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2798:
    begin
        saidaYMax<=352;
        saidaYm<=262;
    end
2799:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2800:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2801:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2802:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2803:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2804:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2805:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2806:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2807:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2808:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2809:
    begin
        saidaYMax<=353;
        saidaYm<=263;
    end
2810:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2811:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2812:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2813:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2814:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2815:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2816:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2817:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2818:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2819:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2820:
    begin
        saidaYMax<=354;
        saidaYm<=264;
    end
2821:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2822:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2823:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2824:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2825:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2826:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2827:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2828:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2829:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2830:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2831:
    begin
        saidaYMax<=355;
        saidaYm<=265;
    end
2832:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2833:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2834:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2835:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2836:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2837:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2838:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2839:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2840:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2841:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2842:
    begin
        saidaYMax<=356;
        saidaYm<=266;
    end
2843:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2844:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2845:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2846:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2847:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2848:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2849:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2850:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2851:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2852:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2853:
    begin
        saidaYMax<=357;
        saidaYm<=267;
    end
2854:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2855:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2856:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2857:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2858:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2859:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2860:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2861:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2862:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2863:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2864:
    begin
        saidaYMax<=358;
        saidaYm<=268;
    end
2865:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2866:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2867:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2868:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2869:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2870:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2871:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2872:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2873:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2874:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2875:
    begin
        saidaYMax<=359;
        saidaYm<=269;
    end
2876:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2877:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2878:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2879:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2880:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2881:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2882:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2883:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2884:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2885:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2886:
    begin
        saidaYMax<=360;
        saidaYm<=270;
    end
2887:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2888:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2889:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2890:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2891:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2892:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2893:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2894:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2895:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2896:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2897:
    begin
        saidaYMax<=361;
        saidaYm<=271;
    end
2898:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2899:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2900:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2901:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2902:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2903:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2904:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2905:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2906:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2907:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2908:
    begin
        saidaYMax<=362;
        saidaYm<=272;
    end
2909:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2910:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2911:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2912:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2913:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2914:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2915:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2916:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2917:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2918:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2919:
    begin
        saidaYMax<=363;
        saidaYm<=273;
    end
2920:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2921:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2922:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2923:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2924:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2925:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2926:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2927:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2928:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2929:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2930:
    begin
        saidaYMax<=364;
        saidaYm<=274;
    end
2931:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2932:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2933:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2934:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2935:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2936:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2937:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2938:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2939:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2940:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2941:
    begin
        saidaYMax<=365;
        saidaYm<=275;
    end
2942:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2943:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2944:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2945:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2946:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2947:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2948:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2949:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2950:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2951:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2952:
    begin
        saidaYMax<=366;
        saidaYm<=276;
    end
2953:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2954:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2955:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2956:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2957:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2958:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2959:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2960:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2961:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2962:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2963:
    begin
        saidaYMax<=367;
        saidaYm<=277;
    end
2964:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2965:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2966:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2967:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2968:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2969:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2970:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2971:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2972:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2973:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2974:
    begin
        saidaYMax<=368;
        saidaYm<=278;
    end
2975:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2976:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2977:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2978:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2979:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2980:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2981:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2982:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2983:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2984:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2985:
    begin
        saidaYMax<=369;
        saidaYm<=279;
    end
2986:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2987:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2988:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2989:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2990:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2991:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2992:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2993:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2994:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2995:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2996:
    begin
        saidaYMax<=370;
        saidaYm<=280;
    end
2997:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
2998:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
2999:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
3000:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
3001:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
3002:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
3003:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
3004:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
3005:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
3006:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
3007:
    begin
        saidaYMax<=371;
        saidaYm<=281;
    end
3008:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3009:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3010:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3011:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3012:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3013:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3014:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3015:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3016:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3017:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3018:
    begin
        saidaYMax<=372;
        saidaYm<=282;
    end
3019:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3020:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3021:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3022:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3023:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3024:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3025:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3026:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3027:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3028:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3029:
    begin
        saidaYMax<=373;
        saidaYm<=283;
    end
3030:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3031:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3032:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3033:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3034:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3035:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3036:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3037:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3038:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3039:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3040:
    begin
        saidaYMax<=374;
        saidaYm<=284;
    end
3041:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3042:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3043:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3044:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3045:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3046:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3047:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3048:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3049:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3050:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3051:
    begin
        saidaYMax<=375;
        saidaYm<=285;
    end
3052:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3053:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3054:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3055:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3056:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3057:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3058:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3059:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3060:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3061:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3062:
    begin
        saidaYMax<=376;
        saidaYm<=286;
    end
3063:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3064:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3065:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3066:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3067:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3068:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3069:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3070:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3071:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3072:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3073:
    begin
        saidaYMax<=377;
        saidaYm<=287;
    end
3074:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3075:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3076:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3077:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3078:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3079:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3080:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3081:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3082:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3083:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3084:
    begin
        saidaYMax<=378;
        saidaYm<=288;
    end
3085:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3086:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3087:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3088:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3089:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3090:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3091:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3092:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3093:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3094:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3095:
    begin
        saidaYMax<=379;
        saidaYm<=289;
    end
3096:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3097:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3098:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3099:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3100:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3101:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3102:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3103:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3104:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3105:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3106:
    begin
        saidaYMax<=380;
        saidaYm<=290;
    end
3107:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3108:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3109:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3110:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3111:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3112:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3113:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3114:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3115:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3116:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3117:
    begin
        saidaYMax<=381;
        saidaYm<=291;
    end
3118:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3119:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3120:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3121:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3122:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3123:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3124:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3125:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3126:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3127:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3128:
    begin
        saidaYMax<=382;
        saidaYm<=292;
    end
3129:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3130:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3131:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3132:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3133:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3134:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3135:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3136:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3137:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3138:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3139:
    begin
        saidaYMax<=383;
        saidaYm<=293;
    end
3140:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3141:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3142:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3143:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3144:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3145:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3146:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3147:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3148:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3149:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3150:
    begin
        saidaYMax<=384;
        saidaYm<=294;
    end
3151:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3152:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3153:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3154:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3155:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3156:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3157:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3158:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3159:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3160:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3161:
    begin
        saidaYMax<=385;
        saidaYm<=295;
    end
3162:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3163:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3164:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3165:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3166:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3167:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3168:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3169:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3170:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3171:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3172:
    begin
        saidaYMax<=386;
        saidaYm<=296;
    end
3173:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3174:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3175:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3176:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3177:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3178:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3179:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3180:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3181:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3182:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3183:
    begin
        saidaYMax<=387;
        saidaYm<=297;
    end
3184:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3185:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3186:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3187:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3188:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3189:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3190:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3191:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3192:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3193:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3194:
    begin
        saidaYMax<=388;
        saidaYm<=298;
    end
3195:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3196:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3197:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3198:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3199:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3200:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3201:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3202:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3203:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3204:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3205:
    begin
        saidaYMax<=389;
        saidaYm<=299;
    end
3206:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3207:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3208:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3209:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3210:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3211:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3212:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3213:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3214:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3215:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3216:
    begin
        saidaYMax<=390;
        saidaYm<=300;
    end
3217:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3218:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3219:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3220:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3221:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3222:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3223:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3224:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3225:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3226:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3227:
    begin
        saidaYMax<=391;
        saidaYm<=301;
    end
3228:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3229:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3230:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3231:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3232:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3233:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3234:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3235:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3236:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3237:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3238:
    begin
        saidaYMax<=392;
        saidaYm<=302;
    end
3239:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3240:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3241:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3242:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3243:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3244:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3245:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3246:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3247:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3248:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3249:
    begin
        saidaYMax<=393;
        saidaYm<=303;
    end
3250:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3251:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3252:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3253:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3254:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3255:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3256:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3257:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3258:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3259:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3260:
    begin
        saidaYMax<=394;
        saidaYm<=304;
    end
3261:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3262:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3263:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3264:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3265:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3266:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3267:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3268:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3269:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3270:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3271:
    begin
        saidaYMax<=395;
        saidaYm<=305;
    end
3272:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3273:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3274:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3275:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3276:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3277:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3278:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3279:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3280:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3281:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3282:
    begin
        saidaYMax<=396;
        saidaYm<=306;
    end
3283:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3284:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3285:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3286:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3287:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3288:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3289:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3290:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3291:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3292:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3293:
    begin
        saidaYMax<=397;
        saidaYm<=307;
    end
3294:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3295:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3296:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3297:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3298:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3299:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3300:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3301:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3302:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3303:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3304:
    begin
        saidaYMax<=398;
        saidaYm<=308;
    end
3305:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3306:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3307:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3308:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3309:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3310:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3311:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3312:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3313:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3314:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3315:
    begin
        saidaYMax<=399;
        saidaYm<=309;
    end
3316:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3317:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3318:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3319:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3320:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3321:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3322:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3323:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3324:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3325:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3326:
    begin
        saidaYMax<=400;
        saidaYm<=310;
    end
3327:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3328:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3329:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3330:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3331:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3332:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3333:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3334:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3335:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3336:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3337:
    begin
        saidaYMax<=401;
        saidaYm<=311;
    end
3338:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3339:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3340:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3341:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3342:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3343:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3344:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3345:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3346:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3347:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3348:
    begin
        saidaYMax<=402;
        saidaYm<=312;
    end
3349:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3350:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3351:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3352:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3353:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3354:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3355:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3356:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3357:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3358:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3359:
    begin
        saidaYMax<=403;
        saidaYm<=313;
    end
3360:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3361:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3362:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3363:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3364:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3365:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3366:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3367:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3368:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3369:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3370:
    begin
        saidaYMax<=404;
        saidaYm<=314;
    end
3371:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3372:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3373:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3374:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3375:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3376:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3377:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3378:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3379:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3380:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3381:
    begin
        saidaYMax<=405;
        saidaYm<=315;
    end
3382:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3383:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3384:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3385:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3386:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3387:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3388:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3389:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3390:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3391:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3392:
    begin
        saidaYMax<=406;
        saidaYm<=316;
    end
3393:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3394:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3395:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3396:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3397:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3398:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3399:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3400:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3401:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3402:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3403:
    begin
        saidaYMax<=407;
        saidaYm<=317;
    end
3404:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3405:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3406:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3407:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3408:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3409:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3410:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3411:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3412:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3413:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3414:
    begin
        saidaYMax<=408;
        saidaYm<=318;
    end
3415:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3416:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3417:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3418:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3419:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3420:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3421:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3422:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3423:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3424:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3425:
    begin
        saidaYMax<=409;
        saidaYm<=319;
    end
3426:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3427:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3428:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3429:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3430:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3431:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3432:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3433:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3434:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3435:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3436:
    begin
        saidaYMax<=410;
        saidaYm<=320;
    end
3437:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3438:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3439:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3440:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3441:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3442:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3443:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3444:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3445:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3446:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3447:
    begin
        saidaYMax<=411;
        saidaYm<=321;
    end
3448:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3449:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3450:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3451:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3452:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3453:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3454:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3455:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3456:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3457:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3458:
    begin
        saidaYMax<=412;
        saidaYm<=322;
    end
3459:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3460:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3461:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3462:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3463:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3464:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3465:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3466:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3467:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3468:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3469:
    begin
        saidaYMax<=413;
        saidaYm<=323;
    end
3470:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3471:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3472:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3473:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3474:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3475:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3476:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3477:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3478:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3479:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3480:
    begin
        saidaYMax<=414;
        saidaYm<=324;
    end
3481:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3482:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3483:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3484:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3485:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3486:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3487:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3488:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3489:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3490:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3491:
    begin
        saidaYMax<=415;
        saidaYm<=325;
    end
3492:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3493:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3494:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3495:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3496:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3497:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3498:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3499:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3500:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3501:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3502:
    begin
        saidaYMax<=416;
        saidaYm<=326;
    end
3503:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3504:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3505:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3506:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3507:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3508:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3509:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3510:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3511:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3512:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3513:
    begin
        saidaYMax<=417;
        saidaYm<=327;
    end
3514:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3515:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3516:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3517:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3518:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3519:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3520:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3521:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3522:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3523:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3524:
    begin
        saidaYMax<=418;
        saidaYm<=328;
    end
3525:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3526:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3527:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3528:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3529:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3530:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3531:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3532:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3533:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3534:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3535:
    begin
        saidaYMax<=419;
        saidaYm<=329;
    end
3536:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3537:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3538:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3539:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3540:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3541:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3542:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3543:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3544:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3545:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3546:
    begin
        saidaYMax<=420;
        saidaYm<=330;
    end
3547:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3548:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3549:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3550:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3551:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3552:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3553:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3554:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3555:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3556:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3557:
    begin
        saidaYMax<=421;
        saidaYm<=331;
    end
3558:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3559:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3560:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3561:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3562:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3563:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3564:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3565:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3566:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3567:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3568:
    begin
        saidaYMax<=422;
        saidaYm<=332;
    end
3569:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3570:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3571:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3572:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3573:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3574:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3575:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3576:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3577:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3578:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3579:
    begin
        saidaYMax<=423;
        saidaYm<=333;
    end
3580:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3581:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3582:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3583:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3584:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3585:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3586:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3587:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3588:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3589:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3590:
    begin
        saidaYMax<=424;
        saidaYm<=334;
    end
3591:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3592:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3593:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3594:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3595:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3596:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3597:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3598:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3599:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3600:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3601:
    begin
        saidaYMax<=425;
        saidaYm<=335;
    end
3602:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3603:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3604:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3605:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3606:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3607:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3608:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3609:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3610:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3611:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3612:
    begin
        saidaYMax<=426;
        saidaYm<=336;
    end
3613:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3614:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3615:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3616:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3617:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3618:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3619:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3620:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3621:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3622:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3623:
    begin
        saidaYMax<=427;
        saidaYm<=337;
    end
3624:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3625:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3626:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3627:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3628:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3629:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3630:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3631:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3632:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3633:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3634:
    begin
        saidaYMax<=428;
        saidaYm<=338;
    end
3635:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3636:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3637:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3638:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3639:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3640:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3641:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3642:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3643:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3644:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3645:
    begin
        saidaYMax<=429;
        saidaYm<=339;
    end
3646:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3647:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3648:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3649:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3650:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3651:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3652:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3653:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3654:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3655:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3656:
    begin
        saidaYMax<=430;
        saidaYm<=340;
    end
3657:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3658:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3659:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3660:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3661:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3662:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3663:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3664:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3665:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3666:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3667:
    begin
        saidaYMax<=431;
        saidaYm<=341;
    end
3668:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3669:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3670:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3671:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3672:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3673:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3674:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3675:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3676:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3677:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3678:
    begin
        saidaYMax<=432;
        saidaYm<=342;
    end
3679:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3680:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3681:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3682:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3683:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3684:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3685:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3686:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3687:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3688:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3689:
    begin
        saidaYMax<=433;
        saidaYm<=343;
    end
3690:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3691:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3692:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3693:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3694:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3695:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3696:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3697:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3698:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3699:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3700:
    begin
        saidaYMax<=434;
        saidaYm<=344;
    end
3701:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3702:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3703:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3704:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3705:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3706:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3707:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3708:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3709:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3710:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3711:
    begin
        saidaYMax<=435;
        saidaYm<=345;
    end
3712:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3713:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3714:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3715:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3716:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3717:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3718:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3719:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3720:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3721:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3722:
    begin
        saidaYMax<=436;
        saidaYm<=346;
    end
3723:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3724:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3725:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3726:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3727:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3728:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3729:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3730:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3731:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3732:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3733:
    begin
        saidaYMax<=437;
        saidaYm<=347;
    end
3734:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3735:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3736:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3737:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3738:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3739:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3740:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3741:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3742:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3743:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3744:
    begin
        saidaYMax<=438;
        saidaYm<=348;
    end
3745:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3746:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3747:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3748:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3749:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3750:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3751:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3752:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3753:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3754:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3755:
    begin
        saidaYMax<=439;
        saidaYm<=349;
    end
3756:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3757:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3758:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3759:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3760:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3761:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3762:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3763:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3764:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3765:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3766:
    begin
        saidaYMax<=440;
        saidaYm<=350;
    end
3767:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3768:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3769:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3770:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3771:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3772:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3773:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3774:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3775:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3776:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3777:
    begin
        saidaYMax<=441;
        saidaYm<=351;
    end
3778:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3779:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3780:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3781:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3782:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3783:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3784:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3785:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3786:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3787:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3788:
    begin
        saidaYMax<=442;
        saidaYm<=352;
    end
3789:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3790:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3791:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3792:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3793:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3794:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3795:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3796:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3797:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3798:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3799:
    begin
        saidaYMax<=443;
        saidaYm<=353;
    end
3800:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3801:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3802:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3803:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3804:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3805:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3806:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3807:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3808:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3809:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3810:
    begin
        saidaYMax<=444;
        saidaYm<=354;
    end
3811:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3812:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3813:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3814:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3815:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3816:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3817:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3818:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3819:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3820:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3821:
    begin
        saidaYMax<=445;
        saidaYm<=355;
    end
3822:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3823:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3824:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3825:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3826:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3827:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3828:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3829:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3830:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3831:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3832:
    begin
        saidaYMax<=446;
        saidaYm<=356;
    end
3833:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3834:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3835:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3836:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3837:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3838:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3839:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3840:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3841:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3842:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3843:
    begin
        saidaYMax<=447;
        saidaYm<=357;
    end
3844:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3845:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3846:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3847:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3848:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3849:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3850:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3851:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3852:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3853:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3854:
    begin
        saidaYMax<=448;
        saidaYm<=358;
    end
3855:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3856:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3857:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3858:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3859:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3860:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3861:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3862:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3863:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3864:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3865:
    begin
        saidaYMax<=449;
        saidaYm<=359;
    end
3866:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3867:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3868:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3869:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3870:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3871:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3872:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3873:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3874:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3875:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3876:
    begin
        saidaYMax<=450;
        saidaYm<=360;
    end
3877:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3878:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3879:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3880:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3881:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3882:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3883:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3884:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3885:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3886:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3887:
    begin
        saidaYMax<=451;
        saidaYm<=361;
    end
3888:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3889:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3890:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3891:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3892:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3893:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3894:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3895:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3896:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3897:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3898:
    begin
        saidaYMax<=452;
        saidaYm<=362;
    end
3899:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3900:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3901:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3902:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3903:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3904:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3905:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3906:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3907:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3908:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3909:
    begin
        saidaYMax<=453;
        saidaYm<=363;
    end
3910:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3911:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3912:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3913:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3914:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3915:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3916:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3917:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3918:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3919:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3920:
    begin
        saidaYMax<=454;
        saidaYm<=364;
    end
3921:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3922:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3923:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3924:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3925:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3926:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3927:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3928:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3929:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3930:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3931:
    begin
        saidaYMax<=455;
        saidaYm<=365;
    end
3932:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3933:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3934:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3935:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3936:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3937:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3938:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3939:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3940:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3941:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3942:
    begin
        saidaYMax<=456;
        saidaYm<=366;
    end
3943:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3944:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3945:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3946:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3947:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3948:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3949:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3950:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3951:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3952:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3953:
    begin
        saidaYMax<=457;
        saidaYm<=367;
    end
3954:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3955:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3956:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3957:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3958:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3959:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3960:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3961:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3962:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3963:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3964:
    begin
        saidaYMax<=458;
        saidaYm<=368;
    end
3965:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3966:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3967:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3968:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3969:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3970:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3971:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3972:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3973:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3974:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3975:
    begin
        saidaYMax<=459;
        saidaYm<=369;
    end
3976:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3977:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3978:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3979:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3980:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3981:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3982:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3983:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3984:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3985:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3986:
    begin
        saidaYMax<=460;
        saidaYm<=370;
    end
3987:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3988:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3989:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3990:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3991:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3992:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3993:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3994:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3995:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3996:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3997:
    begin
        saidaYMax<=461;
        saidaYm<=371;
    end
3998:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
3999:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
4000:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
4001:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
4002:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
4003:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
4004:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
4005:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
4006:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
4007:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
4008:
    begin
        saidaYMax<=462;
        saidaYm<=372;
    end
4009:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4010:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4011:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4012:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4013:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4014:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4015:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4016:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4017:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4018:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4019:
    begin
        saidaYMax<=463;
        saidaYm<=373;
    end
4020:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4021:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4022:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4023:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4024:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4025:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4026:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4027:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4028:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4029:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4030:
    begin
        saidaYMax<=464;
        saidaYm<=374;
    end
4031:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4032:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4033:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4034:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4035:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4036:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4037:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4038:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4039:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4040:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4041:
    begin
        saidaYMax<=465;
        saidaYm<=375;
    end
4042:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4043:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4044:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4045:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4046:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4047:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4048:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4049:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4050:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4051:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4052:
    begin
        saidaYMax<=466;
        saidaYm<=376;
    end
4053:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4054:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4055:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4056:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4057:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4058:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4059:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4060:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4061:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4062:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4063:
    begin
        saidaYMax<=467;
        saidaYm<=377;
    end
4064:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4065:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4066:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4067:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4068:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4069:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4070:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4071:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4072:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4073:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4074:
    begin
        saidaYMax<=468;
        saidaYm<=378;
    end
4075:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4076:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4077:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4078:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4079:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4080:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4081:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4082:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4083:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4084:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4085:
    begin
        saidaYMax<=469;
        saidaYm<=379;
    end
4086:
    begin
        saidaYMax<=470;
        saidaYm<=380;
    end
4087:
    begin
        saidaYMax<=470;
        saidaYm<=380;
    end
4088:
    begin
        saidaYMax<=470;
        saidaYm<=380;
    end
4089:
    begin
        saidaYMax<=470;
        saidaYm<=380;
    end
4090:
    begin
        saidaYMax<=470;
        saidaYm<=380;
    end
4091:
    begin
        saidaYMax<=470;
        saidaYm<=380;
    end
4092:
    begin
        saidaYMax<=470;
        saidaYm<=380;
    end
4093:
    begin
        saidaYMax<=470;
        saidaYm<=380;
    end
4094:
    begin
        saidaYMax<=470;
        saidaYm<=380;
    end
4095:
    begin
        saidaYMax<=470;
        saidaYm<=380;
    end
endcase
end
endmodule
