module Teste(output reg [10:0] palete2aux=95);




endmodule

