module constanteDados(output reg[10:0] Paleta1YMax,Paleta1YMin,Paleta2YMax,Paleta2YMin,BalaXMax,BolaXMin,BolaYMax,BolaYMin);
initial Paleta1YMax=95;
initial Paleta1YMin=5;
initial Paleta2YMax=200;
initial Paleta2YMin=110;
initial BalaXMax=110;
initial BolaXMin=80;
initial BolaYMax=50;
initial BolaYMin=20;


endmodule
